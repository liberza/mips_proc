module controller(input wire[5:0] op,
						input wire[5:0] func,
						input wire zero,
						input wire clock,
						input wire reset,
						output reg[6:0] muxctrl,
						output reg[1:0] memctrl,
						output reg[2:0] aluctrl
						);
	
endmodule
	